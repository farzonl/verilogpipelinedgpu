//Returns sin(INVAL) where INVAL is in the range [-255,255] in 1.8.7 format

module sine_LUT(INVAL,OUTVAL);
input[15:0] INVAL;
output[15:0] OUTVAL;

//Round INVAL to the nearest degree
wire[15:0] INVAL_rounded = (INVAL[15] == 1 && INVAL[7] == 1'b1) ? {INVAL[15:7] - 1'b1,7'b0} : (INVAL[15] == 0 && INVAL[7] == 1'b1) ? {INVAL[15:7] + 1'b1,7'b0} : {INVAL[15:7],7'b0};

assign OUTVAL = (INVAL_rounded == 16'hd300) ? 16'hff80 : 
				(INVAL_rounded == 16'hd380 || INVAL_rounded == 16'hd280) ? 16'hff80 : 
				(INVAL_rounded == 16'hd400 || INVAL_rounded == 16'hd200) ? 16'hff80 : 
				(INVAL_rounded == 16'hd480 || INVAL_rounded == 16'hd180) ? 16'hff80 : 
				(INVAL_rounded == 16'hd500 || INVAL_rounded == 16'hd100) ? 16'hff80 : 
				(INVAL_rounded == 16'hd580 || INVAL_rounded == 16'hd080) ? 16'hff80 : 
				(INVAL_rounded == 16'hd600 || INVAL_rounded == 16'hd000) ? 16'hff81 : 
				(INVAL_rounded == 16'hd680 || INVAL_rounded == 16'hcf80) ? 16'hff81 : 
				(INVAL_rounded == 16'hd700 || INVAL_rounded == 16'hcf00) ? 16'hff81 : 
				(INVAL_rounded == 16'hd780 || INVAL_rounded == 16'hce80) ? 16'hff82 : 
				(INVAL_rounded == 16'hd800 || INVAL_rounded == 16'hce00) ? 16'hff82 : 
				(INVAL_rounded == 16'hd880 || INVAL_rounded == 16'hcd80) ? 16'hff82 : 
				(INVAL_rounded == 16'hd900 || INVAL_rounded == 16'hcd00) ? 16'hff83 : 
				(INVAL_rounded == 16'hd980 || INVAL_rounded == 16'hcc80) ? 16'hff83 : 
				(INVAL_rounded == 16'hda00 || INVAL_rounded == 16'hcc00) ? 16'hff84 : 
				(INVAL_rounded == 16'hda80 || INVAL_rounded == 16'hcb80) ? 16'hff84 : 
				(INVAL_rounded == 16'hdb00 || INVAL_rounded == 16'hcb00) ? 16'hff85 : 
				(INVAL_rounded == 16'hdb80 || INVAL_rounded == 16'hca80) ? 16'hff86 : 
				(INVAL_rounded == 16'hdc00 || INVAL_rounded == 16'hca00) ? 16'hff86 : 
				(INVAL_rounded == 16'hdc80 || INVAL_rounded == 16'hc980) ? 16'hff87 : 
				(INVAL_rounded == 16'hdd00 || INVAL_rounded == 16'hc900) ? 16'hff88 : 
				(INVAL_rounded == 16'hdd80 || INVAL_rounded == 16'hc880) ? 16'hff89 : 
				(INVAL_rounded == 16'hde00 || INVAL_rounded == 16'hc800) ? 16'hff89 : 
				(INVAL_rounded == 16'hde80 || INVAL_rounded == 16'hc780) ? 16'hff8a : 
				(INVAL_rounded == 16'hdf00 || INVAL_rounded == 16'hc700) ? 16'hff8b : 
				(INVAL_rounded == 16'hdf80 || INVAL_rounded == 16'hc680) ? 16'hff8c : 
				(INVAL_rounded == 16'he000 || INVAL_rounded == 16'hc600) ? 16'hff8d : 
				(INVAL_rounded == 16'he080 || INVAL_rounded == 16'hc580) ? 16'hff8e : 
				(INVAL_rounded == 16'he100 || INVAL_rounded == 16'hc500) ? 16'hff8f : 
				(INVAL_rounded == 16'he180 || INVAL_rounded == 16'hc480) ? 16'hff90 : 
				(INVAL_rounded == 16'he200 || INVAL_rounded == 16'hc400) ? 16'hff91 : 
				(INVAL_rounded == 16'he280 || INVAL_rounded == 16'hc380) ? 16'hff92 : 
				(INVAL_rounded == 16'he300 || INVAL_rounded == 16'hc300) ? 16'hff93 : 
				(INVAL_rounded == 16'he380 || INVAL_rounded == 16'hc280) ? 16'hff95 : 
				(INVAL_rounded == 16'he400 || INVAL_rounded == 16'hc200) ? 16'hff96 : 
				(INVAL_rounded == 16'he480 || INVAL_rounded == 16'hc180) ? 16'hff97 : 
				(INVAL_rounded == 16'he500 || INVAL_rounded == 16'hc100) ? 16'hff98 : 
				(INVAL_rounded == 16'he580 || INVAL_rounded == 16'hc080) ? 16'hff9a : 
				(INVAL_rounded == 16'he600 || INVAL_rounded == 16'hc000) ? 16'hff9b : 
				(INVAL_rounded == 16'he680 || INVAL_rounded == 16'hbf80) ? 16'hff9d : 
				(INVAL_rounded == 16'he700 || INVAL_rounded == 16'hbf00) ? 16'hff9e : 
				(INVAL_rounded == 16'he780 || INVAL_rounded == 16'hbe80) ? 16'hff9f : 
				(INVAL_rounded == 16'he800 || INVAL_rounded == 16'hbe00) ? 16'hffa1 : 
				(INVAL_rounded == 16'he880 || INVAL_rounded == 16'hbd80) ? 16'hffa2 : 
				(INVAL_rounded == 16'he900 || INVAL_rounded == 16'hbd00) ? 16'hffa4 : 
				(INVAL_rounded == 16'he980 || INVAL_rounded == 16'hbc80) ? 16'hffa5 : 
				(INVAL_rounded == 16'hea00 || INVAL_rounded == 16'hbc00) ? 16'hffa7 : 
				(INVAL_rounded == 16'hea80 || INVAL_rounded == 16'hbb80) ? 16'hffa9 : 
				(INVAL_rounded == 16'heb00 || INVAL_rounded == 16'hbb00) ? 16'hffaa : 
				(INVAL_rounded == 16'heb80 || INVAL_rounded == 16'hba80) ? 16'hffac : 
				(INVAL_rounded == 16'hec00 || INVAL_rounded == 16'hba00) ? 16'hffae : 
				(INVAL_rounded == 16'hec80 || INVAL_rounded == 16'hb980) ? 16'hffaf : 
				(INVAL_rounded == 16'hed00 || INVAL_rounded == 16'hb900) ? 16'hffb1 : 
				(INVAL_rounded == 16'hed80 || INVAL_rounded == 16'hb880) ? 16'hffb3 : 
				(INVAL_rounded == 16'hee00 || INVAL_rounded == 16'hb800) ? 16'hffb5 : 
				(INVAL_rounded == 16'hee80 || INVAL_rounded == 16'hb780) ? 16'hffb7 : 
				(INVAL_rounded == 16'hef00 || INVAL_rounded == 16'hb700) ? 16'hffb8 : 
				(INVAL_rounded == 16'hef80 || INVAL_rounded == 16'hb680) ? 16'hffba : 
				(INVAL_rounded == 16'hf000 || INVAL_rounded == 16'hb600) ? 16'hffbc : 
				(INVAL_rounded == 16'hf080 || INVAL_rounded == 16'hb580) ? 16'hffbe : 
				(INVAL_rounded == 16'hf100 || INVAL_rounded == 16'hb500) ? 16'hffc0 : 
				(INVAL_rounded == 16'hf180 || INVAL_rounded == 16'hb480) ? 16'hffc2 : 
				(INVAL_rounded == 16'hf200 || INVAL_rounded == 16'hb400) ? 16'hffc4 : 
				(INVAL_rounded == 16'hf280 || INVAL_rounded == 16'hb380) ? 16'hffc6 : 
				(INVAL_rounded == 16'hf300 || INVAL_rounded == 16'hb300) ? 16'hffc8 : 
				(INVAL_rounded == 16'hf380 || INVAL_rounded == 16'hb280) ? 16'hffca : 
				(INVAL_rounded == 16'hf400 || INVAL_rounded == 16'hb200) ? 16'hffcc : 
				(INVAL_rounded == 16'hf480 || INVAL_rounded == 16'hb180) ? 16'hffce : 
				(INVAL_rounded == 16'hf500 || INVAL_rounded == 16'hb100) ? 16'hffd0 : 
				(INVAL_rounded == 16'hf580 || INVAL_rounded == 16'hb080) ? 16'hffd2 : 
				(INVAL_rounded == 16'hf600 || INVAL_rounded == 16'hb000) ? 16'hffd4 : 
				(INVAL_rounded == 16'hf680 || INVAL_rounded == 16'haf80) ? 16'hffd6 : 
				(INVAL_rounded == 16'hf700 || INVAL_rounded == 16'haf00) ? 16'hffd8 : 
				(INVAL_rounded == 16'hf780 || INVAL_rounded == 16'hae80) ? 16'hffdb : 
				(INVAL_rounded == 16'hf800 || INVAL_rounded == 16'hae00) ? 16'hffdd : 
				(INVAL_rounded == 16'hf880 || INVAL_rounded == 16'had80) ? 16'hffdf : 
				(INVAL_rounded == 16'hf900 || INVAL_rounded == 16'had00) ? 16'hffe1 : 
				(INVAL_rounded == 16'hf980 || INVAL_rounded == 16'hac80) ? 16'hffe3 : 
				(INVAL_rounded == 16'hfa00 || INVAL_rounded == 16'hac00) ? 16'hffe5 : 
				(INVAL_rounded == 16'hfa80 || INVAL_rounded == 16'hab80) ? 16'hffe8 : 
				(INVAL_rounded == 16'hfb00 || INVAL_rounded == 16'hab00) ? 16'hffea : 
				(INVAL_rounded == 16'hfb80 || INVAL_rounded == 16'haa80) ? 16'hffec : 
				(INVAL_rounded == 16'hfc00 || INVAL_rounded == 16'haa00) ? 16'hffee : 
				(INVAL_rounded == 16'hfc80 || INVAL_rounded == 16'ha980) ? 16'hfff0 : 
				(INVAL_rounded == 16'hfd00 || INVAL_rounded == 16'ha900) ? 16'hfff3 : 
				(INVAL_rounded == 16'hfd80 || INVAL_rounded == 16'ha880) ? 16'hfff5 : 
				(INVAL_rounded == 16'hfe00 || INVAL_rounded == 16'ha800) ? 16'hfff7 : 
				(INVAL_rounded == 16'hfe80 || INVAL_rounded == 16'ha780) ? 16'hfff9 : 
				(INVAL_rounded == 16'hff00 || INVAL_rounded == 16'ha700) ? 16'hfffc : 
				(INVAL_rounded == 16'hff80 || INVAL_rounded == 16'ha680) ? 16'hfffe : 
				(INVAL_rounded == 16'h0 || INVAL_rounded == 16'h5a00) ? 16'h0 : 
				(INVAL_rounded == 16'h80 || INVAL_rounded == 16'h5980) ? 16'h2 : 
				(INVAL_rounded == 16'h100 || INVAL_rounded == 16'h5900) ? 16'h4 : 
				(INVAL_rounded == 16'h180 || INVAL_rounded == 16'h5880) ? 16'h7 : 
				(INVAL_rounded == 16'h200 || INVAL_rounded == 16'h5800) ? 16'h9 : 
				(INVAL_rounded == 16'h280 || INVAL_rounded == 16'h5780) ? 16'hb : 
				(INVAL_rounded == 16'h300 || INVAL_rounded == 16'h5700) ? 16'hd : 
				(INVAL_rounded == 16'h380 || INVAL_rounded == 16'h5680) ? 16'h10 : 
				(INVAL_rounded == 16'h400 || INVAL_rounded == 16'h5600) ? 16'h12 : 
				(INVAL_rounded == 16'h480 || INVAL_rounded == 16'h5580) ? 16'h14 : 
				(INVAL_rounded == 16'h500 || INVAL_rounded == 16'h5500) ? 16'h16 : 
				(INVAL_rounded == 16'h580 || INVAL_rounded == 16'h5480) ? 16'h18 : 
				(INVAL_rounded == 16'h600 || INVAL_rounded == 16'h5400) ? 16'h1b : 
				(INVAL_rounded == 16'h680 || INVAL_rounded == 16'h5380) ? 16'h1d : 
				(INVAL_rounded == 16'h700 || INVAL_rounded == 16'h5300) ? 16'h1f : 
				(INVAL_rounded == 16'h780 || INVAL_rounded == 16'h5280) ? 16'h21 : 
				(INVAL_rounded == 16'h800 || INVAL_rounded == 16'h5200) ? 16'h23 : 
				(INVAL_rounded == 16'h880 || INVAL_rounded == 16'h5180) ? 16'h25 : 
				(INVAL_rounded == 16'h900 || INVAL_rounded == 16'h5100) ? 16'h28 : 
				(INVAL_rounded == 16'h980 || INVAL_rounded == 16'h5080) ? 16'h2a : 
				(INVAL_rounded == 16'ha00 || INVAL_rounded == 16'h5000) ? 16'h2c : 
				(INVAL_rounded == 16'ha80 || INVAL_rounded == 16'h4f80) ? 16'h2e : 
				(INVAL_rounded == 16'hb00 || INVAL_rounded == 16'h4f00) ? 16'h30 : 
				(INVAL_rounded == 16'hb80 || INVAL_rounded == 16'h4e80) ? 16'h32 : 
				(INVAL_rounded == 16'hc00 || INVAL_rounded == 16'h4e00) ? 16'h34 : 
				(INVAL_rounded == 16'hc80 || INVAL_rounded == 16'h4d80) ? 16'h36 : 
				(INVAL_rounded == 16'hd00 || INVAL_rounded == 16'h4d00) ? 16'h38 : 
				(INVAL_rounded == 16'hd80 || INVAL_rounded == 16'h4c80) ? 16'h3a : 
				(INVAL_rounded == 16'he00 || INVAL_rounded == 16'h4c00) ? 16'h3c : 
				(INVAL_rounded == 16'he80 || INVAL_rounded == 16'h4b80) ? 16'h3e : 
				(INVAL_rounded == 16'hf00 || INVAL_rounded == 16'h4b00) ? 16'h40 : 
				(INVAL_rounded == 16'hf80 || INVAL_rounded == 16'h4a80) ? 16'h42 : 
				(INVAL_rounded == 16'h1000 || INVAL_rounded == 16'h4a00) ? 16'h44 : 
				(INVAL_rounded == 16'h1080 || INVAL_rounded == 16'h4980) ? 16'h46 : 
				(INVAL_rounded == 16'h1100 || INVAL_rounded == 16'h4900) ? 16'h48 : 
				(INVAL_rounded == 16'h1180 || INVAL_rounded == 16'h4880) ? 16'h49 : 
				(INVAL_rounded == 16'h1200 || INVAL_rounded == 16'h4800) ? 16'h4b : 
				(INVAL_rounded == 16'h1280 || INVAL_rounded == 16'h4780) ? 16'h4d : 
				(INVAL_rounded == 16'h1300 || INVAL_rounded == 16'h4700) ? 16'h4f : 
				(INVAL_rounded == 16'h1380 || INVAL_rounded == 16'h4680) ? 16'h51 : 
				(INVAL_rounded == 16'h1400 || INVAL_rounded == 16'h4600) ? 16'h52 : 
				(INVAL_rounded == 16'h1480 || INVAL_rounded == 16'h4580) ? 16'h54 : 
				(INVAL_rounded == 16'h1500 || INVAL_rounded == 16'h4500) ? 16'h56 : 
				(INVAL_rounded == 16'h1580 || INVAL_rounded == 16'h4480) ? 16'h57 : 
				(INVAL_rounded == 16'h1600 || INVAL_rounded == 16'h4400) ? 16'h59 : 
				(INVAL_rounded == 16'h1680 || INVAL_rounded == 16'h4380) ? 16'h5b : 
				(INVAL_rounded == 16'h1700 || INVAL_rounded == 16'h4300) ? 16'h5c : 
				(INVAL_rounded == 16'h1780 || INVAL_rounded == 16'h4280) ? 16'h5e : 
				(INVAL_rounded == 16'h1800 || INVAL_rounded == 16'h4200) ? 16'h5f : 
				(INVAL_rounded == 16'h1880 || INVAL_rounded == 16'h4180) ? 16'h61 : 
				(INVAL_rounded == 16'h1900 || INVAL_rounded == 16'h4100) ? 16'h62 : 
				(INVAL_rounded == 16'h1980 || INVAL_rounded == 16'h4080) ? 16'h63 : 
				(INVAL_rounded == 16'h1a00 || INVAL_rounded == 16'h4000) ? 16'h65 : 
				(INVAL_rounded == 16'h1a80 || INVAL_rounded == 16'h3f80) ? 16'h66 : 
				(INVAL_rounded == 16'h1b00 || INVAL_rounded == 16'h3f00) ? 16'h68 : 
				(INVAL_rounded == 16'h1b80 || INVAL_rounded == 16'h3e80) ? 16'h69 : 
				(INVAL_rounded == 16'h1c00 || INVAL_rounded == 16'h3e00) ? 16'h6a : 
				(INVAL_rounded == 16'h1c80 || INVAL_rounded == 16'h3d80) ? 16'h6b : 
				(INVAL_rounded == 16'h1d00 || INVAL_rounded == 16'h3d00) ? 16'h6d : 
				(INVAL_rounded == 16'h1d80 || INVAL_rounded == 16'h3c80) ? 16'h6e : 
				(INVAL_rounded == 16'h1e00 || INVAL_rounded == 16'h3c00) ? 16'h6f : 
				(INVAL_rounded == 16'h1e80 || INVAL_rounded == 16'h3b80) ? 16'h70 : 
				(INVAL_rounded == 16'h1f00 || INVAL_rounded == 16'h3b00) ? 16'h71 : 
				(INVAL_rounded == 16'h1f80 || INVAL_rounded == 16'h3a80) ? 16'h72 : 
				(INVAL_rounded == 16'h2000 || INVAL_rounded == 16'h3a00) ? 16'h73 : 
				(INVAL_rounded == 16'h2080 || INVAL_rounded == 16'h3980) ? 16'h74 : 
				(INVAL_rounded == 16'h2100 || INVAL_rounded == 16'h3900) ? 16'h75 : 
				(INVAL_rounded == 16'h2180 || INVAL_rounded == 16'h3880) ? 16'h76 : 
				(INVAL_rounded == 16'h2200 || INVAL_rounded == 16'h3800) ? 16'h77 : 
				(INVAL_rounded == 16'h2280 || INVAL_rounded == 16'h3780) ? 16'h77 : 
				(INVAL_rounded == 16'h2300 || INVAL_rounded == 16'h3700) ? 16'h78 : 
				(INVAL_rounded == 16'h2380 || INVAL_rounded == 16'h3680) ? 16'h79 : 
				(INVAL_rounded == 16'h2400 || INVAL_rounded == 16'h3600) ? 16'h7a : 
				(INVAL_rounded == 16'h2480 || INVAL_rounded == 16'h3580) ? 16'h7a : 
				(INVAL_rounded == 16'h2500 || INVAL_rounded == 16'h3500) ? 16'h7b : 
				(INVAL_rounded == 16'h2580 || INVAL_rounded == 16'h3480) ? 16'h7c : 
				(INVAL_rounded == 16'h2600 || INVAL_rounded == 16'h3400) ? 16'h7c : 
				(INVAL_rounded == 16'h2680 || INVAL_rounded == 16'h3380) ? 16'h7d : 
				(INVAL_rounded == 16'h2700 || INVAL_rounded == 16'h3300) ? 16'h7d : 
				(INVAL_rounded == 16'h2780 || INVAL_rounded == 16'h3280) ? 16'h7e : 
				(INVAL_rounded == 16'h2800 || INVAL_rounded == 16'h3200) ? 16'h7e : 
				(INVAL_rounded == 16'h2880 || INVAL_rounded == 16'h3180) ? 16'h7e : 
				(INVAL_rounded == 16'h2900 || INVAL_rounded == 16'h3100) ? 16'h7f : 
				(INVAL_rounded == 16'h2980 || INVAL_rounded == 16'h3080) ? 16'h7f : 
				(INVAL_rounded == 16'h2a00 || INVAL_rounded == 16'h3000) ? 16'h7f : 
				(INVAL_rounded == 16'h2a80 || INVAL_rounded == 16'h2f80) ? 16'h80 : 
				(INVAL_rounded == 16'h2b00 || INVAL_rounded == 16'h2f00) ? 16'h80 : 
				(INVAL_rounded == 16'h2b80 || INVAL_rounded == 16'h2e80) ? 16'h80 : 
				(INVAL_rounded == 16'h2c00 || INVAL_rounded == 16'h2e00) ? 16'h80 : 
				(INVAL_rounded == 16'h2c80 || INVAL_rounded == 16'h2d80) ? 16'h80 : 
				(INVAL_rounded == 16'h2d00) ? 16'h80 : 16'hXXXX;
endmodule
